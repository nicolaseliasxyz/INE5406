library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity somador_8_unsigned is
    port(a, b: in std_logic_vector(7 downto 0);
        s: out std_logic_vector(7 downto 0));

end somador_8_unsigned;

architecture comportamento of somador_8_unsigned is
begin

    s <= a + b;

end comportamento;